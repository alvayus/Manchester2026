
library ieee;
use ieee.std_logic_1164.all;
use work.okt_global_pkg.all;
use work.okt_cu_pkg.all;
use work.okt_imu_pkg.all;

entity okt_cu is                        -- Control Unit
    Port(
        clk       : out   std_logic;    -- 100.8 MHz
        rst_n     : in    std_logic;
        -- USB 3.0 interface
        okUH      : in    std_logic_vector(OK_UH_WIDTH_BUS - 1 downto 0);
        okHU      : out   std_logic_vector(OK_HU_WIDTH_BUS - 1 downto 0);
        okUHU     : inout std_logic_vector(OK_UHU_WIDTH_BUS - 1 downto 0);
        okAA      : inout std_logic;
        -- Data in interface
        ecu_data  : in    std_logic_vector(BUFFER_BITS_WIDTH - 1 downto 0);
        ecu_rd    : out   std_logic;
        ecu_ready : in    std_logic;
        -- Input selection
        input_sel : out   std_logic_vector(NUM_INPUTS - 1 downto 0)
    );
end okt_cu;

architecture Behavioral of okt_cu is

    signal n_command   : std_logic_vector(COMMAND_BIT_WIDTH - 1 downto 0);
    signal n_input_sel : std_logic_vector(NUM_INPUTS - 1 downto 0);

    -- ECU Signals
    signal n_ecu_data  : std_logic_vector(BUFFER_BITS_WIDTH - 1 downto 0);
    signal n_ecu_rd    : std_logic;
    signal n_ecu_ready : std_logic;

    -- USB signals
    signal okClk : std_logic;
    signal okHE  : std_logic_vector(OK_HE_WIDTH_BUS - 1 downto 0);
    signal okEH  : std_logic_vector(OK_EH_WIDTH_BUS - 1 downto 0);
    signal okEHx : std_logic_vector(OK_EH_WIDTH_BUS * OK_NUM_okEHx_END_POINTS - 1 downto 0);

    -- OK Endpoints
    signal ep00wire         : std_logic_vector(BUFFER_BITS_WIDTH - 1 downto 0);
    signal ep01wire         : std_logic_vector(BUFFER_BITS_WIDTH - 1 downto 0);
    signal epA0_datain      : std_logic_vector(BUFFER_BITS_WIDTH - 1 downto 0);
    signal epA0_read        : std_logic;
    signal epA0_blockstrobe : std_logic;
    signal epA0_ready       : std_logic;

begin

    n_ecu_data  <= ecu_data;
    ecu_rd      <= n_ecu_rd;
    n_ecu_ready <= ecu_ready;

    okHI : entity work.okHost
        port map(
            okUH  => okUH,
            okHU  => okHU,
            okUHU => okUHU,
            okAA  => okAA,
            okClk => okClk,             -- 100.8 MHz
            okHE  => okHE,
            okEH  => okEH
        );
    clk <= okClk;

    okOR : entity work.okWireOR
        generic map(
            N => OK_NUM_okEHx_END_POINTS
        )
        port map(
            okEH  => okEH,
            okEHx => okEHx
        );

    cmd_EP : entity work.okWireIn
        port map(
            okHE       => okHE,
            ep_addr    => x"00",
            ep_dataout => ep00wire
        );
    n_command <= ep00wire(COMMAND_BIT_WIDTH - 1 downto 0);

    selInput_EP : entity work.okWireIn
        port map(
            okHE       => okHE,
            ep_addr    => x"01",
            ep_dataout => ep01wire
        );
    n_input_sel <= ep01wire(NUM_INPUTS - 1 downto 0);
    input_sel   <= n_input_sel;

    data_out_EP : entity work.okBTPipeOut
        port map(
            okHE           => okHE,
            okEH           => okEHx(1 * OK_EH_WIDTH_BUS - 1 downto 0 * OK_EH_WIDTH_BUS),
            ep_addr        => x"A0",
            ep_read        => epA0_read,
            ep_blockstrobe => epA0_blockstrobe,
            ep_datain      => epA0_datain,
            ep_ready       => epA0_ready
        );

    command_multiplexer : process(n_command, epA0_read, n_ecu_data, n_ecu_ready)
    begin
        n_ecu_rd    <= '0';
        epA0_datain <= (others => '0');
        epA0_ready  <= '0';

        if (n_command(0) = '1') then    -- Send out captured event to USB
            n_ecu_rd    <= epA0_read;
            epA0_datain <= n_ecu_data;
            epA0_ready  <= n_ecu_ready;
        end if;
    end process;

end Behavioral;

