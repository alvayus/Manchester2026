//------------------------------------------------------------------------
// ramtest.v
//
// This sample uses the Xilinx MIG DDR4 controller and HDL to move data
// from the PC to the DDR4 and vice-versa. Based on MIG generated example_top.v.
//
// Host Interface registers:
// WireIn 0x00
//     0 - DDR4 read enable (0=disabled, 1=enabled)
//     1 - DDR4 write enable (0=disabled, 1=enabled)
//     2 - Reset
//
// PipeIn 0x80 - DDR4 write port (U11, DDR2)
// PipeOut 0xA0 - DDR4 read port (U11, DDR2)
//
// This sample is included for reference only.  No guarantees, either
// expressed or implied, are to be drawn.
//------------------------------------------------------------------------
// tabstop 3
// Copyright (c) 2005-2022 Opal Kelly Incorporated
// $Rev$ $Date$
//------------------------------------------------------------------------
`timescale 1ns/1ps
`default_nettype none

module ramtest (
	input  wire [4:0]   okUH,
	output wire [2:0]   okHU,
	inout  wire [31:0]  okUHU,
	inout  wire         okAA,

	input  wire         ddr4_refclk_p,
	input  wire         ddr4_refclk_n,
	
	output wire [5:0]   led,
	
	inout  wire [15:0]  ddr4_dq,
	inout  wire [1:0]   ddr4_dqs_t,
	inout  wire [1:0]   ddr4_dqs_c,
	inout  wire [1:0]   ddr4_dm,
	output wire [0:0]   ddr4_act_n,
	output wire [16:0]  ddr4_addr,
	output wire [1 :0]  ddr4_ba,
	output wire [0:0]   ddr4_bg,
	output wire [0 :0]  ddr4_ck_t,
	output wire [0 :0]  ddr4_ck_c,
	output wire [0 :0]  ddr4_cke,
	output wire [0 :0]  ddr4_cs_n,
	output wire [0 :0]  ddr4_odt,
	output wire         ddr4_reset_n
	);

// OK RAMTest Parameters
localparam BLOCK_SIZE = 128; // 512 bytes / 4 bytes per word, 
localparam FIFO_SIZE = 1023; // note that Xilinx does not allow use of the full 1024 words
localparam BUFFER_HEADROOM = 20; // headroom for the FIFO count to account for latency

// Capability bitfield, used to indicate features supported by this bitfile:
// [0] - Supports passing calibration status through FrontPanel
localparam CAPABILITY = 16'h0001;


wire          init_calib_complete;
reg           sys_rst;

wire [28 :0]  app_addr;
wire [2  :0]  app_cmd;
wire          app_en;
wire          app_rdy;
wire [127:0]  app_rd_data;
wire          app_rd_data_end;
wire          app_rd_data_valid;
wire [127:0]  app_wdf_data;
wire                       app_wdf_end;
wire [15 :0]  app_wdf_mask;
wire          app_wdf_rdy;
wire          app_wdf_wren;

wire          clk;
wire          rst;

// Front Panel

// Target interface bus:
wire         okClk;
wire [112:0] okHE;
wire [64:0]  okEH;

wire [31:0]  ep00wire;

wire         pipe_in_read;
wire [127:0] pipe_in_data;
wire [7:0]   pipe_in_rd_count;
wire [9:0]   pipe_in_wr_count;
wire         pipe_in_valid;
wire         pipe_in_full;
wire         pipe_in_empty;
reg          pipe_in_ready;

wire         pipe_out_write;
wire [127:0] pipe_out_data;
wire [9:0]   pipe_out_rd_count;
wire [7:0]   pipe_out_wr_count;
wire         pipe_out_full;
wire         pipe_out_empty;
reg          pipe_out_ready;

// Pipe Fifos
wire         pi0_ep_write;
wire         po0_ep_read;
wire [31:0]  pi0_ep_dataout;
wire [31:0]  po0_ep_datain;

assign led = {2'b00, ep00wire[0],ep00wire[1],app_wdf_rdy,init_calib_complete};

	//MIG Infrastructure Reset
reg [31:0] rst_cnt;
initial rst_cnt = 32'b0;
always @(posedge okClk) begin
	if(rst_cnt < 32'h0000_0001) begin // minimum 5 ns reset pulse (PG150)
		rst_cnt <= rst_cnt + 1;		  // 1 okClk cycle is 9.92 ns
		sys_rst <= 1'b1;
	end
	else begin
		sys_rst <= 1'b0;
	end
end

// MIG User Interface instantiation
ddr4_0 ddr4_0_i (
  .c0_init_calib_complete   (init_calib_complete),  // output wire c0_init_calib_complete
  .dbg_clk                  (),                     // output wire dbg_clk
  .c0_sys_clk_p             (ddr4_refclk_p),        // input wire c0_sys_clk_p
  .c0_sys_clk_n             (ddr4_refclk_n),        // input wire c0_sys_clk_n
  .dbg_bus                  (),                     // output wire [511 : 0] dbg_bus
  .c0_ddr4_adr              (ddr4_addr),            // output wire [16 : 0] c0_ddr4_adr
  .c0_ddr4_ba               (ddr4_ba),              // output wire [1 : 0] c0_ddr4_ba
  .c0_ddr4_cke              (ddr4_cke),             // output wire [0 : 0] c0_ddr4_cke
  .c0_ddr4_cs_n             (ddr4_cs_n),            // output wire [0 : 0] c0_ddr4_cs_n
  .c0_ddr4_dm_dbi_n         (ddr4_dm),              // inout wire [1 : 0] c0_ddr4_dm_dbi_n
  .c0_ddr4_dq               (ddr4_dq),              // inout wire [15 : 0] c0_ddr4_dq
  .c0_ddr4_dqs_c            (ddr4_dqs_c),           // inout wire [1 : 0] c0_ddr4_dqs_c
  .c0_ddr4_dqs_t            (ddr4_dqs_t),           // inout wire [1 : 0] c0_ddr4_dqs_t
  .c0_ddr4_odt              (ddr4_odt),             // output wire [0 : 0] c0_ddr4_odt
  .c0_ddr4_bg               (ddr4_bg),              // output wire [0 : 0] c0_ddr4_bg
  .c0_ddr4_reset_n          (ddr4_reset_n),         // output wire c0_ddr4_reset_n
  .c0_ddr4_act_n            (ddr4_act_n),           // output wire c0_ddr4_act_n
  .c0_ddr4_ck_c             (ddr4_ck_c),            // output wire [0 : 0] c0_ddr4_ck_c
  .c0_ddr4_ck_t             (ddr4_ck_t),            // output wire [0 : 0] c0_ddr4_ck_t
  
  .c0_ddr4_ui_clk           (clk),                  // output wire c0_ddr4_ui_clk
  .c0_ddr4_ui_clk_sync_rst  (rst),                  // output wire c0_ddr4_ui_clk_sync_rst
  
  .c0_ddr4_app_en           (app_en),               // input wire c0_ddr4_app_en
  .c0_ddr4_app_hi_pri       (1'b0),                 // input wire c0_ddr4_app_hi_pri
  .c0_ddr4_app_wdf_end      (app_wdf_end),          // input wire c0_ddr4_app_wdf_end
  .c0_ddr4_app_wdf_wren     (app_wdf_wren),         // input wire c0_ddr4_app_wdf_wren
  .c0_ddr4_app_rd_data_end  (app_rd_data_end),      // output wire c0_ddr4_app_rd_data_end
  .c0_ddr4_app_rd_data_valid(app_rd_data_valid),    // output wire c0_ddr4_app_rd_data_valid
  .c0_ddr4_app_rdy          (app_rdy),              // output wire c0_ddr4_app_rdy
  .c0_ddr4_app_wdf_rdy      (app_wdf_rdy),          // output wire c0_ddr4_app_wdf_rdy
  .c0_ddr4_app_addr         (app_addr),             // input wire [28 : 0] c0_ddr4_app_addr
  .c0_ddr4_app_cmd          (app_cmd),              // input wire [2 : 0] c0_ddr4_app_cmd
  .c0_ddr4_app_wdf_data     (app_wdf_data),         // input wire [127 : 0] c0_ddr4_app_wdf_data
  .c0_ddr4_app_wdf_mask     (app_wdf_mask),         // input wire [15 : 0] c0_ddr4_app_wdf_mask
  .c0_ddr4_app_rd_data      (app_rd_data),          // output wire [127 : 0] c0_ddr4_app_rd_data
 
  .sys_rst                  (sys_rst)               // input wire sys_rst
);

// OK MIG DDR3 Testbench Instatiation
ddr4_test ddr4_tb (
	.clk                (clk),
	.reset              (ep00wire[2] | rst),
	.reads_en           (ep00wire[0]),
	.writes_en          (ep00wire[1]),
	.calib_done         (init_calib_complete),

	.ib_re              (pipe_in_read),
	.ib_data            (pipe_in_data),
	.ib_count           (pipe_in_rd_count),
	.ib_valid           (pipe_in_valid),
	.ib_empty           (pipe_in_empty),
	
	.ob_we              (pipe_out_write),
	.ob_data            (pipe_out_data),
	.ob_count           (pipe_out_wr_count),
	.ob_full            (pipe_out_full),
	
	.app_rdy            (app_rdy),
	.app_en             (app_en),
	.app_cmd            (app_cmd),
	.app_addr           (app_addr),
	
	.app_rd_data        (app_rd_data),
	.app_rd_data_end    (app_rd_data_end),
	.app_rd_data_valid  (app_rd_data_valid),
	
	.app_wdf_rdy        (app_wdf_rdy),
	.app_wdf_wren       (app_wdf_wren),
	.app_wdf_data       (app_wdf_data),
	.app_wdf_end        (app_wdf_end),
	.app_wdf_mask       (app_wdf_mask)
	);

//Block Throttle
always @(posedge okClk) begin
	// Check for enough space in input FIFO to pipe in another block
	// The count is compared against a reduced size to account for delays in
	// FIFO count updates.
	if(pipe_in_wr_count <= (FIFO_SIZE-BUFFER_HEADROOM-BLOCK_SIZE) ) begin
		pipe_in_ready <= 1'b1;
	end
	else begin
		pipe_in_ready <= 1'b0;
	end

	// Check for enough space in output FIFO to pipe out another block
	if(pipe_out_rd_count >= BLOCK_SIZE) begin
		pipe_out_ready <= 1'b1;
	end
	else begin
		pipe_out_ready <= 1'b0;
	end
end


// Instantiate the okHost and connect endpoints.
wire [65*4-1:0]  okEHx;

okHost okHI(
	.okUH(okUH),
	.okHU(okHU),
	.okUHU(okUHU),
	.okAA(okAA),
	.okClk(okClk),
	.okHE(okHE),
	.okEH(okEH)
	);

okWireOR # (.N(4)) wireOR (okEH, okEHx);
okWireIn       wi00 (.okHE(okHE),                             .ep_addr(8'h00), .ep_dataout(ep00wire));
okWireOut      wo00 (.okHE(okHE), .okEH(okEHx[ 0*65 +: 65 ]), .ep_addr(8'h20), .ep_datain({31'h00, init_calib_complete}));
okWireOut      wo01 (.okHE(okHE), .okEH(okEHx[ 1*65 +: 65 ]), .ep_addr(8'h3e), .ep_datain(CAPABILITY));
okBTPipeIn     pi0  (.okHE(okHE), .okEH(okEHx[ 2*65 +: 65 ]), .ep_addr(8'h80), .ep_write(pi0_ep_write), .ep_blockstrobe(), .ep_dataout(pi0_ep_dataout), .ep_ready(pipe_in_ready));
okBTPipeOut    po0  (.okHE(okHE), .okEH(okEHx[ 3*65 +: 65 ]), .ep_addr(8'ha0), .ep_read(po0_ep_read),   .ep_blockstrobe(), .ep_datain(po0_ep_datain),   .ep_ready(pipe_out_ready));

fifo_w32_1024_r128_256 okPipeIn_fifo (
  .rst          (ep00wire[2]),       // input wire rst
  .wr_clk       (okClk),             // input wire wr_clk
  .rd_clk       (clk),               // input wire rd_clk
  .din          (pi0_ep_dataout),    // input wire [31 : 0] din
  .wr_en        (pi0_ep_write),      // input wire wr_en
  .rd_en        (pipe_in_read),      // input wire rd_en
  .dout         (pipe_in_data),      // output wire [127 : 0] dout
  .full         (pipe_in_full),      // output wire full
  .empty        (pipe_in_empty),     // output wire empty
  .valid        (pipe_in_valid),     // output wire valid
  .rd_data_count(pipe_in_rd_count),  // output wire [7 : 0] rd_data_count
  .wr_data_count(pipe_in_wr_count),  // output wire [9 : 0] wr_data_count
  .wr_rst_busy  (),                  // output wire wr_rst_busy
  .rd_rst_busy  ()                   // output wire rd_rst_busy
);

fifo_w128_256_r32_1024 okPipeOut_fifo (
  .rst          (ep00wire[2]),       // input wire rst
  .wr_clk       (clk),               // input wire wr_clk
  .rd_clk       (okClk),             // input wire rd_clk
  .din          (pipe_out_data),     // input wire [127 : 0] din
  .wr_en        (pipe_out_write),    // input wire wr_en
  .rd_en        (po0_ep_read),       // input wire rd_en
  .dout         (po0_ep_datain),     // output wire [31 : 0] dout
  .full         (pipe_out_full),     // output wire full
  .empty        (pipe_out_empty),    // output wire empty
  .valid        (),                  // output wire valid
  .rd_data_count(pipe_out_rd_count), // output wire [9 : 0] rd_data_count
  .wr_data_count(pipe_out_wr_count), // output wire [7 : 0] wr_data_count
  .wr_rst_busy  (),                  // output wire wr_rst_busy
  .rd_rst_busy  ()                   // output wire rd_rst_busy
);
endmodule
`default_nettype wire
