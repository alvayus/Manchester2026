
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package okt_top_pkg is
	constant ROME_DATA_BITS_WIDTH      : integer := 16;
	constant NODE_DATA_BITS_WIDTH      : integer := 28;
	constant SPINNAKER_BITS_DATA_WIDTH : integer := 8;
end okt_top_pkg;

package body okt_top_pkg is

end okt_top_pkg;
