library ieee;
use ieee.std_logic_1164.all;
use work.okt_global_pkg.all;

package okt_cu_pkg is
    --constant COMMAND_BIT_WIDTH : integer := 3; -- ECU, PASSTROUGH
    --	constant MODE_BUS_WIDTH		: integer := 4;
end okt_cu_pkg;

package body okt_cu_pkg is

end okt_cu_pkg;
