library ieee;
use ieee.STD_LOGIC_1164.all;

package okt_fifo_pkg is
    constant FIFO_ALM_FULL_OFFSET : integer := 64; --before: 64
	 constant FIFO_ALM_EMPTY_OFFSET : integer := 1024; --before: 64
end okt_fifo_pkg;

package body okt_fifo_pkg is
end okt_fifo_pkg;
