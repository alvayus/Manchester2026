library ieee;
use ieee.STD_LOGIC_1164.all;

package okt_fifo_pkg is
<<<<<<< HEAD
    constant FIFO_ALM_FULL_OFFSET : integer := 64; --before: 64
	 constant FIFO_ALM_EMPTY_OFFSET : integer := 64; --before: 64
=======
    constant FIFO_ALM_FULL_OFFSET : integer := 256; --before: 64
	 constant FIFO_ALM_EMPTY_OFFSET : integer := 256; --before: 64
>>>>>>> c0ea32db7e0068b5c23ff21752dd02823d580492
end okt_fifo_pkg;

package body okt_fifo_pkg is
end okt_fifo_pkg;
